// Written by the Majesty Logic Package
module top (
			a[0] , a[1] , a[2] , a[3] , a[4] , a[5] , a[6] , a[7] , a[8] , a[9] , a[10] , a[11] , a[12] , a[13] , a[14] , a[15] , a[16] , a[17] , a[18] , a[19] , a[20] , a[21] , a[22] , a[23] , a[24] , a[25] , a[26] , a[27] , a[28] , a[29] , a[30] , a[31] , a[32] , a[33] , a[34] , a[35] , a[36] , a[37] , a[38] , a[39] , a[40] , a[41] , a[42] , a[43] , a[44] , a[45] , a[46] , a[47] , a[48] , a[49] , a[50] , a[51] , a[52] , a[53] , a[54] , a[55] , a[56] , a[57] , a[58] , a[59] , a[60] , a[61] , a[62] , a[63] , a[64] , a[65] , a[66] , a[67] , a[68] , a[69] , a[70] , a[71] , a[72] , a[73] , a[74] , a[75] , a[76] , a[77] , a[78] , a[79] , a[80] , a[81] , a[82] , a[83] , a[84] , a[85] , a[86] , a[87] , a[88] , a[89] , a[90] , a[91] , a[92] , a[93] , a[94] , a[95] , a[96] , a[97] , a[98] , a[99] , a[100] , a[101] , a[102] , a[103] , a[104] , a[105] , a[106] , a[107] , a[108] , a[109] , a[110] , a[111] , a[112] , a[113] , a[114] , a[115] , a[116] , a[117] , a[118] , a[119] , a[120] , a[121] , a[122] , a[123] , a[124] , a[125] , a[126] , a[127] , b[0] , b[1] , b[2] , b[3] , b[4] , b[5] , b[6] , b[7] , b[8] , b[9] , b[10] , b[11] , b[12] , b[13] , b[14] , b[15] , b[16] , b[17] , b[18] , b[19] , b[20] , b[21] , b[22] , b[23] , b[24] , b[25] , b[26] , b[27] , b[28] , b[29] , b[30] , b[31] , b[32] , b[33] , b[34] , b[35] , b[36] , b[37] , b[38] , b[39] , b[40] , b[41] , b[42] , b[43] , b[44] , b[45] , b[46] , b[47] , b[48] , b[49] , b[50] , b[51] , b[52] , b[53] , b[54] , b[55] , b[56] , b[57] , b[58] , b[59] , b[60] , b[61] , b[62] , b[63] , b[64] , b[65] , b[66] , b[67] , b[68] , b[69] , b[70] , b[71] , b[72] , b[73] , b[74] , b[75] , b[76] , b[77] , b[78] , b[79] , b[80] , b[81] , b[82] , b[83] , b[84] , b[85] , b[86] , b[87] , b[88] , b[89] , b[90] , b[91] , b[92] , b[93] , b[94] , b[95] , b[96] , b[97] , b[98] , b[99] , b[100] , b[101] , b[102] , b[103] , b[104] , b[105] , b[106] , b[107] , b[108] , b[109] , b[110] , b[111] , b[112] , b[113] , b[114] , b[115] , b[116] , b[117] , b[118] , b[119] , b[120] , b[121] , b[122] , b[123] , b[124] , b[125] , b[126] , b[127] , 
			f[0] , f[1] , f[2] , f[3] , f[4] , f[5] , f[6] , f[7] , f[8] , f[9] , f[10] , f[11] , f[12] , f[13] , f[14] , f[15] , f[16] , f[17] , f[18] , f[19] , f[20] , f[21] , f[22] , f[23] , f[24] , f[25] , f[26] , f[27] , f[28] , f[29] , f[30] , f[31] , f[32] , f[33] , f[34] , f[35] , f[36] , f[37] , f[38] , f[39] , f[40] , f[41] , f[42] , f[43] , f[44] , f[45] , f[46] , f[47] , f[48] , f[49] , f[50] , f[51] , f[52] , f[53] , f[54] , f[55] , f[56] , f[57] , f[58] , f[59] , f[60] , f[61] , f[62] , f[63] , f[64] , f[65] , f[66] , f[67] , f[68] , f[69] , f[70] , f[71] , f[72] , f[73] , f[74] , f[75] , f[76] , f[77] , f[78] , f[79] , f[80] , f[81] , f[82] , f[83] , f[84] , f[85] , f[86] , f[87] , f[88] , f[89] , f[90] , f[91] , f[92] , f[93] , f[94] , f[95] , f[96] , f[97] , f[98] , f[99] , f[100] , f[101] , f[102] , f[103] , f[104] , f[105] , f[106] , f[107] , f[108] , f[109] , f[110] , f[111] , f[112] , f[113] , f[114] , f[115] , f[116] , f[117] , f[118] , f[119] , f[120] , f[121] , f[122] , f[123] , f[124] , f[125] , f[126] , f[127] , cOut ) ;
input a[0] , a[1] , a[2] , a[3] , a[4] , a[5] , a[6] , a[7] , a[8] , a[9] , a[10] , a[11] , a[12] , a[13] , a[14] , a[15] , a[16] , a[17] , a[18] , a[19] , a[20] , a[21] , a[22] , a[23] , a[24] , a[25] , a[26] , a[27] , a[28] , a[29] , a[30] , a[31] , a[32] , a[33] , a[34] , a[35] , a[36] , a[37] , a[38] , a[39] , a[40] , a[41] , a[42] , a[43] , a[44] , a[45] , a[46] , a[47] , a[48] , a[49] , a[50] , a[51] , a[52] , a[53] , a[54] , a[55] , a[56] , a[57] , a[58] , a[59] , a[60] , a[61] , a[62] , a[63] , a[64] , a[65] , a[66] , a[67] , a[68] , a[69] , a[70] , a[71] , a[72] , a[73] , a[74] , a[75] , a[76] , a[77] , a[78] , a[79] , a[80] , a[81] , a[82] , a[83] , a[84] , a[85] , a[86] , a[87] , a[88] , a[89] , a[90] , a[91] , a[92] , a[93] , a[94] , a[95] , a[96] , a[97] , a[98] , a[99] , a[100] , a[101] , a[102] , a[103] , a[104] , a[105] , a[106] , a[107] , a[108] , a[109] , a[110] , a[111] , a[112] , a[113] , a[114] , a[115] , a[116] , a[117] , a[118] , a[119] , a[120] , a[121] , a[122] , a[123] , a[124] , a[125] , a[126] , a[127] , b[0] , b[1] , b[2] , b[3] , b[4] , b[5] , b[6] , b[7] , b[8] , b[9] , b[10] , b[11] , b[12] , b[13] , b[14] , b[15] , b[16] , b[17] , b[18] , b[19] , b[20] , b[21] , b[22] , b[23] , b[24] , b[25] , b[26] , b[27] , b[28] , b[29] , b[30] , b[31] , b[32] , b[33] , b[34] , b[35] , b[36] , b[37] , b[38] , b[39] , b[40] , b[41] , b[42] , b[43] , b[44] , b[45] , b[46] , b[47] , b[48] , b[49] , b[50] , b[51] , b[52] , b[53] , b[54] , b[55] , b[56] , b[57] , b[58] , b[59] , b[60] , b[61] , b[62] , b[63] , b[64] , b[65] , b[66] , b[67] , b[68] , b[69] , b[70] , b[71] , b[72] , b[73] , b[74] , b[75] , b[76] , b[77] , b[78] , b[79] , b[80] , b[81] , b[82] , b[83] , b[84] , b[85] , b[86] , b[87] , b[88] , b[89] , b[90] , b[91] , b[92] , b[93] , b[94] , b[95] , b[96] , b[97] , b[98] , b[99] , b[100] , b[101] , b[102] , b[103] , b[104] , b[105] , b[106] , b[107] , b[108] , b[109] , b[110] , b[111] , b[112] , b[113] , b[114] , b[115] , b[116] , b[117] , b[118] , b[119] , b[120] , b[121] , b[122] , b[123] , b[124] , b[125] , b[126] , b[127] ;
output f[0] , f[1] , f[2] , f[3] , f[4] , f[5] , f[6] , f[7] , f[8] , f[9] , f[10] , f[11] , f[12] , f[13] , f[14] , f[15] , f[16] , f[17] , f[18] , f[19] , f[20] , f[21] , f[22] , f[23] , f[24] , f[25] , f[26] , f[27] , f[28] , f[29] , f[30] , f[31] , f[32] , f[33] , f[34] , f[35] , f[36] , f[37] , f[38] , f[39] , f[40] , f[41] , f[42] , f[43] , f[44] , f[45] , f[46] , f[47] , f[48] , f[49] , f[50] , f[51] , f[52] , f[53] , f[54] , f[55] , f[56] , f[57] , f[58] , f[59] , f[60] , f[61] , f[62] , f[63] , f[64] , f[65] , f[66] , f[67] , f[68] , f[69] , f[70] , f[71] , f[72] , f[73] , f[74] , f[75] , f[76] , f[77] , f[78] , f[79] , f[80] , f[81] , f[82] , f[83] , f[84] , f[85] , f[86] , f[87] , f[88] , f[89] , f[90] , f[91] , f[92] , f[93] , f[94] , f[95] , f[96] , f[97] , f[98] , f[99] , f[100] , f[101] , f[102] , f[103] , f[104] , f[105] , f[106] , f[107] , f[108] , f[109] , f[110] , f[111] , f[112] , f[113] , f[114] , f[115] , f[116] , f[117] , f[118] , f[119] , f[120] , f[121] , f[122] , f[123] , f[124] , f[125] , f[126] , f[127] , cOut ;
wire w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 ;
assign w257 = ~a[0] | b[0] ;
assign w258 = a[0] | ~b[0] ;
assign w259 = a[0] & b[0] ;
assign w260 = a[1] | b[1] ;
assign w261 = a[1] & b[1] ;
assign w262 = a[2] | b[2] ;
assign w263 = a[2] & b[2] ;
assign w264 = a[3] | b[3] ;
assign w265 = a[3] & b[3] ;
assign w266 = a[4] | b[4] ;
assign w267 = a[4] & b[4] ;
assign w268 = a[5] | b[5] ;
assign w269 = a[5] & b[5] ;
assign w270 = a[6] | b[6] ;
assign w271 = a[6] & b[6] ;
assign w272 = a[7] | b[7] ;
assign w273 = a[7] & b[7] ;
assign w274 = a[8] | b[8] ;
assign w275 = a[8] & b[8] ;
assign w276 = a[9] | b[9] ;
assign w277 = a[9] & b[9] ;
assign w278 = a[10] | b[10] ;
assign w279 = a[10] & b[10] ;
assign w280 = a[11] | b[11] ;
assign w281 = a[11] & b[11] ;
assign w282 = a[12] | b[12] ;
assign w283 = a[12] & b[12] ;
assign w284 = a[13] | b[13] ;
assign w285 = a[13] & b[13] ;
assign w286 = a[14] | b[14] ;
assign w287 = a[14] & b[14] ;
assign w288 = a[15] | b[15] ;
assign w289 = a[15] & b[15] ;
assign w290 = a[16] | b[16] ;
assign w291 = a[16] & b[16] ;
assign w292 = a[17] | b[17] ;
assign w293 = a[17] & b[17] ;
assign w294 = a[18] | b[18] ;
assign w295 = a[18] & b[18] ;
assign w296 = a[19] | b[19] ;
assign w297 = a[19] & b[19] ;
assign w298 = a[20] | b[20] ;
assign w299 = a[20] & b[20] ;
assign w300 = a[21] | b[21] ;
assign w301 = a[21] & b[21] ;
assign w302 = a[22] | b[22] ;
assign w303 = a[22] & b[22] ;
assign w304 = a[23] | b[23] ;
assign w305 = a[23] & b[23] ;
assign w306 = a[24] | b[24] ;
assign w307 = a[24] & b[24] ;
assign w308 = a[25] | b[25] ;
assign w309 = a[25] & b[25] ;
assign w310 = a[26] | b[26] ;
assign w311 = a[26] & b[26] ;
assign w312 = a[27] | b[27] ;
assign w313 = a[27] & b[27] ;
assign w314 = a[28] | b[28] ;
assign w315 = a[28] & b[28] ;
assign w316 = a[29] | b[29] ;
assign w317 = a[29] & b[29] ;
assign w318 = a[30] | b[30] ;
assign w319 = a[30] & b[30] ;
assign w320 = a[31] | b[31] ;
assign w321 = a[31] & b[31] ;
assign w322 = a[32] | b[32] ;
assign w323 = a[32] & b[32] ;
assign w324 = a[33] | b[33] ;
assign w325 = a[33] & b[33] ;
assign w326 = a[34] | b[34] ;
assign w327 = a[34] & b[34] ;
assign w328 = a[35] | b[35] ;
assign w329 = a[35] & b[35] ;
assign w330 = a[36] | b[36] ;
assign w331 = a[36] & b[36] ;
assign w332 = a[37] | b[37] ;
assign w333 = a[37] & b[37] ;
assign w334 = a[38] | b[38] ;
assign w335 = a[38] & b[38] ;
assign w336 = a[39] | b[39] ;
assign w337 = a[39] & b[39] ;
assign w338 = a[40] | b[40] ;
assign w339 = a[40] & b[40] ;
assign w340 = a[41] | b[41] ;
assign w341 = a[41] & b[41] ;
assign w342 = a[42] | b[42] ;
assign w343 = a[42] & b[42] ;
assign w344 = a[43] | b[43] ;
assign w345 = a[43] & b[43] ;
assign w346 = a[44] | b[44] ;
assign w347 = a[44] & b[44] ;
assign w348 = a[45] | b[45] ;
assign w349 = a[45] & b[45] ;
assign w350 = a[46] | b[46] ;
assign w351 = a[46] & b[46] ;
assign w352 = a[47] | b[47] ;
assign w353 = a[47] & b[47] ;
assign w354 = a[48] | b[48] ;
assign w355 = a[48] & b[48] ;
assign w356 = a[49] | b[49] ;
assign w357 = a[49] & b[49] ;
assign w358 = a[50] | b[50] ;
assign w359 = a[50] & b[50] ;
assign w360 = a[51] | b[51] ;
assign w361 = a[51] & b[51] ;
assign w362 = a[52] | b[52] ;
assign w363 = a[52] & b[52] ;
assign w364 = a[53] | b[53] ;
assign w365 = a[53] & b[53] ;
assign w366 = a[54] | b[54] ;
assign w367 = a[54] & b[54] ;
assign w368 = a[55] | b[55] ;
assign w369 = a[55] & b[55] ;
assign w370 = a[56] | b[56] ;
assign w371 = a[56] & b[56] ;
assign w372 = a[57] | b[57] ;
assign w373 = a[57] & b[57] ;
assign w374 = a[58] | b[58] ;
assign w375 = a[58] & b[58] ;
assign w376 = a[59] | b[59] ;
assign w377 = a[59] & b[59] ;
assign w378 = a[60] | b[60] ;
assign w379 = a[60] & b[60] ;
assign w380 = a[61] | b[61] ;
assign w381 = a[61] & b[61] ;
assign w382 = a[62] | b[62] ;
assign w383 = a[62] & b[62] ;
assign w384 = a[63] | b[63] ;
assign w385 = a[63] & b[63] ;
assign w386 = a[64] | b[64] ;
assign w387 = a[64] & b[64] ;
assign w388 = a[65] | b[65] ;
assign w389 = a[65] & b[65] ;
assign w390 = a[66] | b[66] ;
assign w391 = a[66] & b[66] ;
assign w392 = a[67] | b[67] ;
assign w393 = a[67] & b[67] ;
assign w394 = a[68] | b[68] ;
assign w395 = a[68] & b[68] ;
assign w396 = a[69] | b[69] ;
assign w397 = a[69] & b[69] ;
assign w398 = a[70] | b[70] ;
assign w399 = a[70] & b[70] ;
assign w400 = a[71] | b[71] ;
assign w401 = a[71] & b[71] ;
assign w402 = a[72] | b[72] ;
assign w403 = a[72] & b[72] ;
assign w404 = a[73] | b[73] ;
assign w405 = a[73] & b[73] ;
assign w406 = a[74] | b[74] ;
assign w407 = a[74] & b[74] ;
assign w408 = a[75] | b[75] ;
assign w409 = a[75] & b[75] ;
assign w410 = a[76] | b[76] ;
assign w411 = a[76] & b[76] ;
assign w412 = a[77] | b[77] ;
assign w413 = a[77] & b[77] ;
assign w414 = a[78] | b[78] ;
assign w415 = a[78] & b[78] ;
assign w416 = a[79] | b[79] ;
assign w417 = a[79] & b[79] ;
assign w418 = a[80] | b[80] ;
assign w419 = a[80] & b[80] ;
assign w420 = a[81] | b[81] ;
assign w421 = a[81] & b[81] ;
assign w422 = a[82] | b[82] ;
assign w423 = a[82] & b[82] ;
assign w424 = a[83] | b[83] ;
assign w425 = a[83] & b[83] ;
assign w426 = a[84] | b[84] ;
assign w427 = a[84] & b[84] ;
assign w428 = a[85] | b[85] ;
assign w429 = a[85] & b[85] ;
assign w430 = a[86] | b[86] ;
assign w431 = a[86] & b[86] ;
assign w432 = a[87] | b[87] ;
assign w433 = a[87] & b[87] ;
assign w434 = a[88] | b[88] ;
assign w435 = a[88] & b[88] ;
assign w436 = a[89] | b[89] ;
assign w437 = a[89] & b[89] ;
assign w438 = a[90] | b[90] ;
assign w439 = a[90] & b[90] ;
assign w440 = a[91] | b[91] ;
assign w441 = a[91] & b[91] ;
assign w442 = a[92] | b[92] ;
assign w443 = a[92] & b[92] ;
assign w444 = a[93] | b[93] ;
assign w445 = a[93] & b[93] ;
assign w446 = a[94] | b[94] ;
assign w447 = a[94] & b[94] ;
assign w448 = a[95] | b[95] ;
assign w449 = a[95] & b[95] ;
assign w450 = a[96] | b[96] ;
assign w451 = a[96] & b[96] ;
assign w452 = a[97] | b[97] ;
assign w453 = a[97] & b[97] ;
assign w454 = a[98] | b[98] ;
assign w455 = a[98] & b[98] ;
assign w456 = a[99] | b[99] ;
assign w457 = a[99] & b[99] ;
assign w458 = a[100] | b[100] ;
assign w459 = a[100] & b[100] ;
assign w460 = a[101] | b[101] ;
assign w461 = a[101] & b[101] ;
assign w462 = a[102] | b[102] ;
assign w463 = a[102] & b[102] ;
assign w464 = a[103] | b[103] ;
assign w465 = a[103] & b[103] ;
assign w466 = a[104] | b[104] ;
assign w467 = a[104] & b[104] ;
assign w468 = a[105] | b[105] ;
assign w469 = a[105] & b[105] ;
assign w470 = a[106] | b[106] ;
assign w471 = a[106] & b[106] ;
assign w472 = a[107] | b[107] ;
assign w473 = a[107] & b[107] ;
assign w474 = a[108] | b[108] ;
assign w475 = a[108] & b[108] ;
assign w476 = a[109] | b[109] ;
assign w477 = a[109] & b[109] ;
assign w478 = a[110] | b[110] ;
assign w479 = a[110] & b[110] ;
assign w480 = a[111] | b[111] ;
assign w481 = a[111] & b[111] ;
assign w482 = a[112] | b[112] ;
assign w483 = a[112] & b[112] ;
assign w484 = a[113] | b[113] ;
assign w485 = a[113] & b[113] ;
assign w486 = a[114] | b[114] ;
assign w487 = a[114] & b[114] ;
assign w488 = a[115] | b[115] ;
assign w489 = a[115] & b[115] ;
assign w490 = a[116] | b[116] ;
assign w491 = a[116] & b[116] ;
assign w492 = a[117] | b[117] ;
assign w493 = a[117] & b[117] ;
assign w494 = a[118] | b[118] ;
assign w495 = a[118] & b[118] ;
assign w496 = a[119] | b[119] ;
assign w497 = a[119] & b[119] ;
assign w498 = a[120] | b[120] ;
assign w499 = a[120] & b[120] ;
assign w500 = a[121] | b[121] ;
assign w501 = a[121] & b[121] ;
assign w502 = a[122] | b[122] ;
assign w503 = a[122] & b[122] ;
assign w504 = a[123] | b[123] ;
assign w505 = a[123] & b[123] ;
assign w506 = a[124] | b[124] ;
assign w507 = a[124] & b[124] ;
assign w508 = a[125] | b[125] ;
assign w509 = a[125] & b[125] ;
assign w510 = a[126] | b[126] ;
assign w511 = a[126] & b[126] ;
assign w512 = a[127] | b[127] ;
assign w513 = a[127] & b[127] ;
assign w514 = w257 & w258 ;
assign w515 = w259 & w260 ;
assign w516 = ~w260 | w261 ;
assign w517 = ~w262 | w263 ;
assign w518 = ~w264 | w265 ;
assign w519 = ~w266 | w267 ;
assign w520 = ~w268 | w269 ;
assign w521 = ~w270 | w271 ;
assign w522 = ~w272 | w273 ;
assign w523 = ~w274 | w275 ;
assign w524 = ~w276 | w277 ;
assign w525 = ~w278 | w279 ;
assign w526 = ~w280 | w281 ;
assign w527 = ~w282 | w283 ;
assign w528 = ~w284 | w285 ;
assign w529 = ~w286 | w287 ;
assign w530 = ~w288 | w289 ;
assign w531 = ~w290 | w291 ;
assign w532 = ~w292 | w293 ;
assign w533 = ~w294 | w295 ;
assign w534 = ~w296 | w297 ;
assign w535 = ~w298 | w299 ;
assign w536 = ~w300 | w301 ;
assign w537 = ~w302 | w303 ;
assign w538 = ~w304 | w305 ;
assign w539 = ~w306 | w307 ;
assign w540 = ~w308 | w309 ;
assign w541 = ~w310 | w311 ;
assign w542 = ~w312 | w313 ;
assign w543 = ~w314 | w315 ;
assign w544 = ~w316 | w317 ;
assign w545 = ~w318 | w319 ;
assign w546 = ~w320 | w321 ;
assign w547 = ~w322 | w323 ;
assign w548 = ~w324 | w325 ;
assign w549 = ~w326 | w327 ;
assign w550 = ~w328 | w329 ;
assign w551 = ~w330 | w331 ;
assign w552 = ~w332 | w333 ;
assign w553 = ~w334 | w335 ;
assign w554 = ~w336 | w337 ;
assign w555 = ~w338 | w339 ;
assign w556 = ~w340 | w341 ;
assign w557 = ~w342 | w343 ;
assign w558 = ~w344 | w345 ;
assign w559 = ~w346 | w347 ;
assign w560 = ~w348 | w349 ;
assign w561 = ~w350 | w351 ;
assign w562 = ~w352 | w353 ;
assign w563 = ~w354 | w355 ;
assign w564 = ~w356 | w357 ;
assign w565 = ~w358 | w359 ;
assign w566 = ~w360 | w361 ;
assign w567 = ~w362 | w363 ;
assign w568 = ~w364 | w365 ;
assign w569 = ~w366 | w367 ;
assign w570 = ~w368 | w369 ;
assign w571 = ~w370 | w371 ;
assign w572 = ~w372 | w373 ;
assign w573 = ~w374 | w375 ;
assign w574 = ~w376 | w377 ;
assign w575 = ~w378 | w379 ;
assign w576 = ~w380 | w381 ;
assign w577 = ~w382 | w383 ;
assign w578 = ~w384 | w385 ;
assign w579 = ~w386 | w387 ;
assign w580 = ~w388 | w389 ;
assign w581 = ~w390 | w391 ;
assign w582 = ~w392 | w393 ;
assign w583 = ~w394 | w395 ;
assign w584 = ~w396 | w397 ;
assign w585 = ~w398 | w399 ;
assign w586 = ~w400 | w401 ;
assign w587 = ~w402 | w403 ;
assign w588 = ~w404 | w405 ;
assign w589 = ~w406 | w407 ;
assign w590 = ~w408 | w409 ;
assign w591 = ~w410 | w411 ;
assign w592 = ~w412 | w413 ;
assign w593 = ~w414 | w415 ;
assign w594 = ~w416 | w417 ;
assign w595 = ~w418 | w419 ;
assign w596 = ~w420 | w421 ;
assign w597 = ~w422 | w423 ;
assign w598 = ~w424 | w425 ;
assign w599 = ~w426 | w427 ;
assign w600 = ~w428 | w429 ;
assign w601 = ~w430 | w431 ;
assign w602 = ~w432 | w433 ;
assign w603 = ~w434 | w435 ;
assign w604 = ~w436 | w437 ;
assign w605 = ~w438 | w439 ;
assign w606 = ~w440 | w441 ;
assign w607 = ~w442 | w443 ;
assign w608 = ~w444 | w445 ;
assign w609 = ~w446 | w447 ;
assign w610 = ~w448 | w449 ;
assign w611 = ~w450 | w451 ;
assign w612 = ~w452 | w453 ;
assign w613 = ~w454 | w455 ;
assign w614 = ~w456 | w457 ;
assign w615 = ~w458 | w459 ;
assign w616 = ~w460 | w461 ;
assign w617 = ~w462 | w463 ;
assign w618 = ~w464 | w465 ;
assign w619 = ~w466 | w467 ;
assign w620 = ~w468 | w469 ;
assign w621 = ~w470 | w471 ;
assign w622 = ~w472 | w473 ;
assign w623 = ~w474 | w475 ;
assign w624 = ~w476 | w477 ;
assign w625 = ~w478 | w479 ;
assign w626 = ~w480 | w481 ;
assign w627 = ~w482 | w483 ;
assign w628 = ~w484 | w485 ;
assign w629 = ~w486 | w487 ;
assign w630 = ~w488 | w489 ;
assign w631 = ~w490 | w491 ;
assign w632 = ~w492 | w493 ;
assign w633 = ~w494 | w495 ;
assign w634 = ~w496 | w497 ;
assign w635 = ~w498 | w499 ;
assign w636 = ~w500 | w501 ;
assign w637 = ~w502 | w503 ;
assign w638 = ~w504 | w505 ;
assign w639 = ~w506 | w507 ;
assign w640 = ~w508 | w509 ;
assign w641 = ~w510 | w511 ;
assign w642 = ~w512 | w513 ;
assign w643 = w261 | w515 ;
assign w644 = w259 & w516 ;
assign w645 = w259 | w516 ;
assign w646 = ~w517 | w643 ;
assign w647 = w517 | ~w643 ;
assign w648 = w262 & w643 ;
assign w649 = w644 | ~w645 ;
assign w650 = w646 & w647 ;
assign w651 = w263 | w648 ;
assign w652 = ~w518 | w651 ;
assign w653 = w518 | ~w651 ;
assign w654 = w264 & w651 ;
assign w655 = w652 & w653 ;
assign w656 = w265 | w654 ;
assign w657 = ~w519 | w656 ;
assign w658 = w519 | ~w656 ;
assign w659 = w266 & w656 ;
assign w660 = w657 & w658 ;
assign w661 = w267 | w659 ;
assign w662 = ~w520 | w661 ;
assign w663 = w520 | ~w661 ;
assign w664 = w268 & w661 ;
assign w665 = w662 & w663 ;
assign w666 = w269 | w664 ;
assign w667 = ~w521 | w666 ;
assign w668 = w521 | ~w666 ;
assign w669 = w270 & w666 ;
assign w670 = w667 & w668 ;
assign w671 = w271 | w669 ;
assign w672 = ~w522 | w671 ;
assign w673 = w522 | ~w671 ;
assign w674 = w272 & w671 ;
assign w675 = w672 & w673 ;
assign w676 = w273 | w674 ;
assign w677 = ~w523 | w676 ;
assign w678 = w523 | ~w676 ;
assign w679 = w274 & w676 ;
assign w680 = w677 & w678 ;
assign w681 = w275 | w679 ;
assign w682 = ~w524 | w681 ;
assign w683 = w524 | ~w681 ;
assign w684 = w276 & w681 ;
assign w685 = w682 & w683 ;
assign w686 = w277 | w684 ;
assign w687 = ~w525 | w686 ;
assign w688 = w525 | ~w686 ;
assign w689 = w278 & w686 ;
assign w690 = w687 & w688 ;
assign w691 = w279 | w689 ;
assign w692 = ~w526 | w691 ;
assign w693 = w526 | ~w691 ;
assign w694 = w280 & w691 ;
assign w695 = w692 & w693 ;
assign w696 = w281 | w694 ;
assign w697 = ~w527 | w696 ;
assign w698 = w527 | ~w696 ;
assign w699 = w282 & w696 ;
assign w700 = w697 & w698 ;
assign w701 = w283 | w699 ;
assign w702 = ~w528 | w701 ;
assign w703 = w528 | ~w701 ;
assign w704 = w284 & w701 ;
assign w705 = w702 & w703 ;
assign w706 = w285 | w704 ;
assign w707 = ~w529 | w706 ;
assign w708 = w529 | ~w706 ;
assign w709 = w286 & w706 ;
assign w710 = w707 & w708 ;
assign w711 = w287 | w709 ;
assign w712 = ~w530 | w711 ;
assign w713 = w530 | ~w711 ;
assign w714 = w288 & w711 ;
assign w715 = w712 & w713 ;
assign w716 = w289 | w714 ;
assign w717 = ~w531 | w716 ;
assign w718 = w531 | ~w716 ;
assign w719 = w290 & w716 ;
assign w720 = w717 & w718 ;
assign w721 = w291 | w719 ;
assign w722 = ~w532 | w721 ;
assign w723 = w532 | ~w721 ;
assign w724 = w292 & w721 ;
assign w725 = w722 & w723 ;
assign w726 = w293 | w724 ;
assign w727 = ~w533 | w726 ;
assign w728 = w533 | ~w726 ;
assign w729 = w294 & w726 ;
assign w730 = w727 & w728 ;
assign w731 = w295 | w729 ;
assign w732 = ~w534 | w731 ;
assign w733 = w534 | ~w731 ;
assign w734 = w296 & w731 ;
assign w735 = w732 & w733 ;
assign w736 = w297 | w734 ;
assign w737 = ~w535 | w736 ;
assign w738 = w535 | ~w736 ;
assign w739 = w298 & w736 ;
assign w740 = w737 & w738 ;
assign w741 = w299 | w739 ;
assign w742 = ~w536 | w741 ;
assign w743 = w536 | ~w741 ;
assign w744 = w300 & w741 ;
assign w745 = w742 & w743 ;
assign w746 = w301 | w744 ;
assign w747 = ~w537 | w746 ;
assign w748 = w537 | ~w746 ;
assign w749 = w302 & w746 ;
assign w750 = w747 & w748 ;
assign w751 = w303 | w749 ;
assign w752 = ~w538 | w751 ;
assign w753 = w538 | ~w751 ;
assign w754 = w304 & w751 ;
assign w755 = w752 & w753 ;
assign w756 = w305 | w754 ;
assign w757 = ~w539 | w756 ;
assign w758 = w539 | ~w756 ;
assign w759 = w306 & w756 ;
assign w760 = w757 & w758 ;
assign w761 = w307 | w759 ;
assign w762 = ~w540 | w761 ;
assign w763 = w540 | ~w761 ;
assign w764 = w308 & w761 ;
assign w765 = w762 & w763 ;
assign w766 = w309 | w764 ;
assign w767 = ~w541 | w766 ;
assign w768 = w541 | ~w766 ;
assign w769 = w310 & w766 ;
assign w770 = w767 & w768 ;
assign w771 = w311 | w769 ;
assign w772 = ~w542 | w771 ;
assign w773 = w542 | ~w771 ;
assign w774 = w312 & w771 ;
assign w775 = w772 & w773 ;
assign w776 = w313 | w774 ;
assign w777 = ~w543 | w776 ;
assign w778 = w543 | ~w776 ;
assign w779 = w314 & w776 ;
assign w780 = w777 & w778 ;
assign w781 = w315 | w779 ;
assign w782 = ~w544 | w781 ;
assign w783 = w544 | ~w781 ;
assign w784 = w316 & w781 ;
assign w785 = w782 & w783 ;
assign w786 = w317 | w784 ;
assign w787 = ~w545 | w786 ;
assign w788 = w545 | ~w786 ;
assign w789 = w318 & w786 ;
assign w790 = w787 & w788 ;
assign w791 = w319 | w789 ;
assign w792 = ~w546 | w791 ;
assign w793 = w546 | ~w791 ;
assign w794 = w320 & w791 ;
assign w795 = w792 & w793 ;
assign w796 = w321 | w794 ;
assign w797 = ~w547 | w796 ;
assign w798 = w547 | ~w796 ;
assign w799 = w322 & w796 ;
assign w800 = w797 & w798 ;
assign w801 = w323 | w799 ;
assign w802 = ~w548 | w801 ;
assign w803 = w548 | ~w801 ;
assign w804 = w324 & w801 ;
assign w805 = w802 & w803 ;
assign w806 = w325 | w804 ;
assign w807 = ~w549 | w806 ;
assign w808 = w549 | ~w806 ;
assign w809 = w326 & w806 ;
assign w810 = w807 & w808 ;
assign w811 = w327 | w809 ;
assign w812 = ~w550 | w811 ;
assign w813 = w550 | ~w811 ;
assign w814 = w328 & w811 ;
assign w815 = w812 & w813 ;
assign w816 = w329 | w814 ;
assign w817 = ~w551 | w816 ;
assign w818 = w551 | ~w816 ;
assign w819 = w330 & w816 ;
assign w820 = w817 & w818 ;
assign w821 = w331 | w819 ;
assign w822 = ~w552 | w821 ;
assign w823 = w552 | ~w821 ;
assign w824 = w332 & w821 ;
assign w825 = w822 & w823 ;
assign w826 = w333 | w824 ;
assign w827 = ~w553 | w826 ;
assign w828 = w553 | ~w826 ;
assign w829 = w334 & w826 ;
assign w830 = w827 & w828 ;
assign w831 = w335 | w829 ;
assign w832 = ~w554 | w831 ;
assign w833 = w554 | ~w831 ;
assign w834 = w336 & w831 ;
assign w835 = w832 & w833 ;
assign w836 = w337 | w834 ;
assign w837 = ~w555 | w836 ;
assign w838 = w555 | ~w836 ;
assign w839 = w338 & w836 ;
assign w840 = w837 & w838 ;
assign w841 = w339 | w839 ;
assign w842 = ~w556 | w841 ;
assign w843 = w556 | ~w841 ;
assign w844 = w340 & w841 ;
assign w845 = w842 & w843 ;
assign w846 = w341 | w844 ;
assign w847 = ~w557 | w846 ;
assign w848 = w557 | ~w846 ;
assign w849 = w342 & w846 ;
assign w850 = w847 & w848 ;
assign w851 = w343 | w849 ;
assign w852 = ~w558 | w851 ;
assign w853 = w558 | ~w851 ;
assign w854 = w344 & w851 ;
assign w855 = w852 & w853 ;
assign w856 = w345 | w854 ;
assign w857 = ~w559 | w856 ;
assign w858 = w559 | ~w856 ;
assign w859 = w346 & w856 ;
assign w860 = w857 & w858 ;
assign w861 = w347 | w859 ;
assign w862 = ~w560 | w861 ;
assign w863 = w560 | ~w861 ;
assign w864 = w348 & w861 ;
assign w865 = w862 & w863 ;
assign w866 = w349 | w864 ;
assign w867 = ~w561 | w866 ;
assign w868 = w561 | ~w866 ;
assign w869 = w350 & w866 ;
assign w870 = w867 & w868 ;
assign w871 = w351 | w869 ;
assign w872 = ~w562 | w871 ;
assign w873 = w562 | ~w871 ;
assign w874 = w352 & w871 ;
assign w875 = w872 & w873 ;
assign w876 = w353 | w874 ;
assign w877 = ~w563 | w876 ;
assign w878 = w563 | ~w876 ;
assign w879 = w354 & w876 ;
assign w880 = w877 & w878 ;
assign w881 = w355 | w879 ;
assign w882 = ~w564 | w881 ;
assign w883 = w564 | ~w881 ;
assign w884 = w356 & w881 ;
assign w885 = w882 & w883 ;
assign w886 = w357 | w884 ;
assign w887 = ~w565 | w886 ;
assign w888 = w565 | ~w886 ;
assign w889 = w358 & w886 ;
assign w890 = w887 & w888 ;
assign w891 = w359 | w889 ;
assign w892 = ~w566 | w891 ;
assign w893 = w566 | ~w891 ;
assign w894 = w360 & w891 ;
assign w895 = w892 & w893 ;
assign w896 = w361 | w894 ;
assign w897 = ~w567 | w896 ;
assign w898 = w567 | ~w896 ;
assign w899 = w362 & w896 ;
assign w900 = w897 & w898 ;
assign w901 = w363 | w899 ;
assign w902 = ~w568 | w901 ;
assign w903 = w568 | ~w901 ;
assign w904 = w364 & w901 ;
assign w905 = w902 & w903 ;
assign w906 = w365 | w904 ;
assign w907 = ~w569 | w906 ;
assign w908 = w569 | ~w906 ;
assign w909 = w366 & w906 ;
assign w910 = w907 & w908 ;
assign w911 = w367 | w909 ;
assign w912 = ~w570 | w911 ;
assign w913 = w570 | ~w911 ;
assign w914 = w368 & w911 ;
assign w915 = w912 & w913 ;
assign w916 = w369 | w914 ;
assign w917 = ~w571 | w916 ;
assign w918 = w571 | ~w916 ;
assign w919 = w370 & w916 ;
assign w920 = w917 & w918 ;
assign w921 = w371 | w919 ;
assign w922 = ~w572 | w921 ;
assign w923 = w572 | ~w921 ;
assign w924 = w372 & w921 ;
assign w925 = w922 & w923 ;
assign w926 = w373 | w924 ;
assign w927 = ~w573 | w926 ;
assign w928 = w573 | ~w926 ;
assign w929 = w374 & w926 ;
assign w930 = w927 & w928 ;
assign w931 = w375 | w929 ;
assign w932 = ~w574 | w931 ;
assign w933 = w574 | ~w931 ;
assign w934 = w376 & w931 ;
assign w935 = w932 & w933 ;
assign w936 = w377 | w934 ;
assign w937 = ~w575 | w936 ;
assign w938 = w575 | ~w936 ;
assign w939 = w378 & w936 ;
assign w940 = w937 & w938 ;
assign w941 = w379 | w939 ;
assign w942 = ~w576 | w941 ;
assign w943 = w576 | ~w941 ;
assign w944 = w380 & w941 ;
assign w945 = w942 & w943 ;
assign w946 = w381 | w944 ;
assign w947 = ~w577 | w946 ;
assign w948 = w577 | ~w946 ;
assign w949 = w382 & w946 ;
assign w950 = w947 & w948 ;
assign w951 = w383 | w949 ;
assign w952 = ~w578 | w951 ;
assign w953 = w578 | ~w951 ;
assign w954 = w384 & w951 ;
assign w955 = w952 & w953 ;
assign w956 = w385 | w954 ;
assign w957 = ~w579 | w956 ;
assign w958 = w579 | ~w956 ;
assign w959 = w386 & w956 ;
assign w960 = w957 & w958 ;
assign w961 = w387 | w959 ;
assign w962 = ~w580 | w961 ;
assign w963 = w580 | ~w961 ;
assign w964 = w388 & w961 ;
assign w965 = w962 & w963 ;
assign w966 = w389 | w964 ;
assign w967 = ~w581 | w966 ;
assign w968 = w581 | ~w966 ;
assign w969 = w390 & w966 ;
assign w970 = w967 & w968 ;
assign w971 = w391 | w969 ;
assign w972 = ~w582 | w971 ;
assign w973 = w582 | ~w971 ;
assign w974 = w392 & w971 ;
assign w975 = w972 & w973 ;
assign w976 = w393 | w974 ;
assign w977 = ~w583 | w976 ;
assign w978 = w583 | ~w976 ;
assign w979 = w394 & w976 ;
assign w980 = w977 & w978 ;
assign w981 = w395 | w979 ;
assign w982 = ~w584 | w981 ;
assign w983 = w584 | ~w981 ;
assign w984 = w396 & w981 ;
assign w985 = w982 & w983 ;
assign w986 = w397 | w984 ;
assign w987 = ~w585 | w986 ;
assign w988 = w585 | ~w986 ;
assign w989 = w398 & w986 ;
assign w990 = w987 & w988 ;
assign w991 = w399 | w989 ;
assign w992 = ~w586 | w991 ;
assign w993 = w586 | ~w991 ;
assign w994 = w400 & w991 ;
assign w995 = w992 & w993 ;
assign w996 = w401 | w994 ;
assign w997 = ~w587 | w996 ;
assign w998 = w587 | ~w996 ;
assign w999 = w402 & w996 ;
assign w1000 = w997 & w998 ;
assign w1001 = w403 | w999 ;
assign w1002 = ~w588 | w1001 ;
assign w1003 = w588 | ~w1001 ;
assign w1004 = w404 & w1001 ;
assign w1005 = w1002 & w1003 ;
assign w1006 = w405 | w1004 ;
assign w1007 = ~w589 | w1006 ;
assign w1008 = w589 | ~w1006 ;
assign w1009 = w406 & w1006 ;
assign w1010 = w1007 & w1008 ;
assign w1011 = w407 | w1009 ;
assign w1012 = ~w590 | w1011 ;
assign w1013 = w590 | ~w1011 ;
assign w1014 = w408 & w1011 ;
assign w1015 = w1012 & w1013 ;
assign w1016 = w409 | w1014 ;
assign w1017 = ~w591 | w1016 ;
assign w1018 = w591 | ~w1016 ;
assign w1019 = w410 & w1016 ;
assign w1020 = w1017 & w1018 ;
assign w1021 = w411 | w1019 ;
assign w1022 = ~w592 | w1021 ;
assign w1023 = w592 | ~w1021 ;
assign w1024 = w412 & w1021 ;
assign w1025 = w1022 & w1023 ;
assign w1026 = w413 | w1024 ;
assign w1027 = ~w593 | w1026 ;
assign w1028 = w593 | ~w1026 ;
assign w1029 = w414 & w1026 ;
assign w1030 = w1027 & w1028 ;
assign w1031 = w415 | w1029 ;
assign w1032 = ~w594 | w1031 ;
assign w1033 = w594 | ~w1031 ;
assign w1034 = w416 & w1031 ;
assign w1035 = w1032 & w1033 ;
assign w1036 = w417 | w1034 ;
assign w1037 = ~w595 | w1036 ;
assign w1038 = w595 | ~w1036 ;
assign w1039 = w418 & w1036 ;
assign w1040 = w1037 & w1038 ;
assign w1041 = w419 | w1039 ;
assign w1042 = ~w596 | w1041 ;
assign w1043 = w596 | ~w1041 ;
assign w1044 = w420 & w1041 ;
assign w1045 = w1042 & w1043 ;
assign w1046 = w421 | w1044 ;
assign w1047 = ~w597 | w1046 ;
assign w1048 = w597 | ~w1046 ;
assign w1049 = w422 & w1046 ;
assign w1050 = w1047 & w1048 ;
assign w1051 = w423 | w1049 ;
assign w1052 = ~w598 | w1051 ;
assign w1053 = w598 | ~w1051 ;
assign w1054 = w424 & w1051 ;
assign w1055 = w1052 & w1053 ;
assign w1056 = w425 | w1054 ;
assign w1057 = ~w599 | w1056 ;
assign w1058 = w599 | ~w1056 ;
assign w1059 = w426 & w1056 ;
assign w1060 = w1057 & w1058 ;
assign w1061 = w427 | w1059 ;
assign w1062 = ~w600 | w1061 ;
assign w1063 = w600 | ~w1061 ;
assign w1064 = w428 & w1061 ;
assign w1065 = w1062 & w1063 ;
assign w1066 = w429 | w1064 ;
assign w1067 = ~w601 | w1066 ;
assign w1068 = w601 | ~w1066 ;
assign w1069 = w430 & w1066 ;
assign w1070 = w1067 & w1068 ;
assign w1071 = w431 | w1069 ;
assign w1072 = ~w602 | w1071 ;
assign w1073 = w602 | ~w1071 ;
assign w1074 = w432 & w1071 ;
assign w1075 = w1072 & w1073 ;
assign w1076 = w433 | w1074 ;
assign w1077 = ~w603 | w1076 ;
assign w1078 = w603 | ~w1076 ;
assign w1079 = w434 & w1076 ;
assign w1080 = w1077 & w1078 ;
assign w1081 = w435 | w1079 ;
assign w1082 = ~w604 | w1081 ;
assign w1083 = w604 | ~w1081 ;
assign w1084 = w436 & w1081 ;
assign w1085 = w1082 & w1083 ;
assign w1086 = w437 | w1084 ;
assign w1087 = ~w605 | w1086 ;
assign w1088 = w605 | ~w1086 ;
assign w1089 = w438 & w1086 ;
assign w1090 = w1087 & w1088 ;
assign w1091 = w439 | w1089 ;
assign w1092 = ~w606 | w1091 ;
assign w1093 = w606 | ~w1091 ;
assign w1094 = w440 & w1091 ;
assign w1095 = w1092 & w1093 ;
assign w1096 = w441 | w1094 ;
assign w1097 = ~w607 | w1096 ;
assign w1098 = w607 | ~w1096 ;
assign w1099 = w442 & w1096 ;
assign w1100 = w1097 & w1098 ;
assign w1101 = w443 | w1099 ;
assign w1102 = ~w608 | w1101 ;
assign w1103 = w608 | ~w1101 ;
assign w1104 = w444 & w1101 ;
assign w1105 = w1102 & w1103 ;
assign w1106 = w445 | w1104 ;
assign w1107 = ~w609 | w1106 ;
assign w1108 = w609 | ~w1106 ;
assign w1109 = w446 & w1106 ;
assign w1110 = w1107 & w1108 ;
assign w1111 = w447 | w1109 ;
assign w1112 = ~w610 | w1111 ;
assign w1113 = w610 | ~w1111 ;
assign w1114 = w448 & w1111 ;
assign w1115 = w1112 & w1113 ;
assign w1116 = w449 | w1114 ;
assign w1117 = ~w611 | w1116 ;
assign w1118 = w611 | ~w1116 ;
assign w1119 = w450 & w1116 ;
assign w1120 = w1117 & w1118 ;
assign w1121 = w451 | w1119 ;
assign w1122 = ~w612 | w1121 ;
assign w1123 = w612 | ~w1121 ;
assign w1124 = w452 & w1121 ;
assign w1125 = w1122 & w1123 ;
assign w1126 = w453 | w1124 ;
assign w1127 = ~w613 | w1126 ;
assign w1128 = w613 | ~w1126 ;
assign w1129 = w454 & w1126 ;
assign w1130 = w1127 & w1128 ;
assign w1131 = w455 | w1129 ;
assign w1132 = ~w614 | w1131 ;
assign w1133 = w614 | ~w1131 ;
assign w1134 = w456 & w1131 ;
assign w1135 = w1132 & w1133 ;
assign w1136 = w457 | w1134 ;
assign w1137 = ~w615 | w1136 ;
assign w1138 = w615 | ~w1136 ;
assign w1139 = w458 & w1136 ;
assign w1140 = w1137 & w1138 ;
assign w1141 = w459 | w1139 ;
assign w1142 = ~w616 | w1141 ;
assign w1143 = w616 | ~w1141 ;
assign w1144 = w460 & w1141 ;
assign w1145 = w1142 & w1143 ;
assign w1146 = w461 | w1144 ;
assign w1147 = ~w617 | w1146 ;
assign w1148 = w617 | ~w1146 ;
assign w1149 = w462 & w1146 ;
assign w1150 = w1147 & w1148 ;
assign w1151 = w463 | w1149 ;
assign w1152 = ~w618 | w1151 ;
assign w1153 = w618 | ~w1151 ;
assign w1154 = w464 & w1151 ;
assign w1155 = w1152 & w1153 ;
assign w1156 = w465 | w1154 ;
assign w1157 = ~w619 | w1156 ;
assign w1158 = w619 | ~w1156 ;
assign w1159 = w466 & w1156 ;
assign w1160 = w1157 & w1158 ;
assign w1161 = w467 | w1159 ;
assign w1162 = ~w620 | w1161 ;
assign w1163 = w620 | ~w1161 ;
assign w1164 = w468 & w1161 ;
assign w1165 = w1162 & w1163 ;
assign w1166 = w469 | w1164 ;
assign w1167 = ~w621 | w1166 ;
assign w1168 = w621 | ~w1166 ;
assign w1169 = w470 & w1166 ;
assign w1170 = w1167 & w1168 ;
assign w1171 = w471 | w1169 ;
assign w1172 = ~w622 | w1171 ;
assign w1173 = w622 | ~w1171 ;
assign w1174 = w472 & w1171 ;
assign w1175 = w1172 & w1173 ;
assign w1176 = w473 | w1174 ;
assign w1177 = ~w623 | w1176 ;
assign w1178 = w623 | ~w1176 ;
assign w1179 = w474 & w1176 ;
assign w1180 = w1177 & w1178 ;
assign w1181 = w475 | w1179 ;
assign w1182 = ~w624 | w1181 ;
assign w1183 = w624 | ~w1181 ;
assign w1184 = w476 & w1181 ;
assign w1185 = w1182 & w1183 ;
assign w1186 = w477 | w1184 ;
assign w1187 = ~w625 | w1186 ;
assign w1188 = w625 | ~w1186 ;
assign w1189 = w478 & w1186 ;
assign w1190 = w1187 & w1188 ;
assign w1191 = w479 | w1189 ;
assign w1192 = ~w626 | w1191 ;
assign w1193 = w626 | ~w1191 ;
assign w1194 = w480 & w1191 ;
assign w1195 = w1192 & w1193 ;
assign w1196 = w481 | w1194 ;
assign w1197 = ~w627 | w1196 ;
assign w1198 = w627 | ~w1196 ;
assign w1199 = w482 & w1196 ;
assign w1200 = w1197 & w1198 ;
assign w1201 = w483 | w1199 ;
assign w1202 = ~w628 | w1201 ;
assign w1203 = w628 | ~w1201 ;
assign w1204 = w484 & w1201 ;
assign w1205 = w1202 & w1203 ;
assign w1206 = w485 | w1204 ;
assign w1207 = ~w629 | w1206 ;
assign w1208 = w629 | ~w1206 ;
assign w1209 = w486 & w1206 ;
assign w1210 = w1207 & w1208 ;
assign w1211 = w487 | w1209 ;
assign w1212 = ~w630 | w1211 ;
assign w1213 = w630 | ~w1211 ;
assign w1214 = w488 & w1211 ;
assign w1215 = w1212 & w1213 ;
assign w1216 = w489 | w1214 ;
assign w1217 = ~w631 | w1216 ;
assign w1218 = w631 | ~w1216 ;
assign w1219 = w490 & w1216 ;
assign w1220 = w1217 & w1218 ;
assign w1221 = w491 | w1219 ;
assign w1222 = ~w632 | w1221 ;
assign w1223 = w632 | ~w1221 ;
assign w1224 = w492 & w1221 ;
assign w1225 = w1222 & w1223 ;
assign w1226 = w493 | w1224 ;
assign w1227 = ~w633 | w1226 ;
assign w1228 = w633 | ~w1226 ;
assign w1229 = w494 & w1226 ;
assign w1230 = w1227 & w1228 ;
assign w1231 = w495 | w1229 ;
assign w1232 = ~w634 | w1231 ;
assign w1233 = w634 | ~w1231 ;
assign w1234 = w496 & w1231 ;
assign w1235 = w1232 & w1233 ;
assign w1236 = w497 | w1234 ;
assign w1237 = ~w635 | w1236 ;
assign w1238 = w635 | ~w1236 ;
assign w1239 = w498 & w1236 ;
assign w1240 = w1237 & w1238 ;
assign w1241 = w499 | w1239 ;
assign w1242 = ~w636 | w1241 ;
assign w1243 = w636 | ~w1241 ;
assign w1244 = w500 & w1241 ;
assign w1245 = w1242 & w1243 ;
assign w1246 = w501 | w1244 ;
assign w1247 = ~w637 | w1246 ;
assign w1248 = w637 | ~w1246 ;
assign w1249 = w502 & w1246 ;
assign w1250 = w1247 & w1248 ;
assign w1251 = w503 | w1249 ;
assign w1252 = ~w638 | w1251 ;
assign w1253 = w638 | ~w1251 ;
assign w1254 = w504 & w1251 ;
assign w1255 = w1252 & w1253 ;
assign w1256 = w505 | w1254 ;
assign w1257 = ~w639 | w1256 ;
assign w1258 = w639 | ~w1256 ;
assign w1259 = w506 & w1256 ;
assign w1260 = w1257 & w1258 ;
assign w1261 = w507 | w1259 ;
assign w1262 = ~w640 | w1261 ;
assign w1263 = w640 | ~w1261 ;
assign w1264 = w508 & w1261 ;
assign w1265 = w1262 & w1263 ;
assign w1266 = w509 | w1264 ;
assign w1267 = ~w641 | w1266 ;
assign w1268 = w641 | ~w1266 ;
assign w1269 = w510 & w1266 ;
assign w1270 = w1267 & w1268 ;
assign w1271 = w511 | w1269 ;
assign w1272 = ~w642 | w1271 ;
assign w1273 = w642 | ~w1271 ;
assign w1274 = w512 & w1271 ;
assign w1275 = w1272 & w1273 ;
assign w1276 = w513 | w1274 ;
assign f[0] = ~w514 ;
assign f[1] = w649 ;
assign f[2] = w650 ;
assign f[3] = w655 ;
assign f[4] = w660 ;
assign f[5] = w665 ;
assign f[6] = w670 ;
assign f[7] = w675 ;
assign f[8] = w680 ;
assign f[9] = w685 ;
assign f[10] = w690 ;
assign f[11] = w695 ;
assign f[12] = w700 ;
assign f[13] = w705 ;
assign f[14] = w710 ;
assign f[15] = w715 ;
assign f[16] = w720 ;
assign f[17] = w725 ;
assign f[18] = w730 ;
assign f[19] = w735 ;
assign f[20] = w740 ;
assign f[21] = w745 ;
assign f[22] = w750 ;
assign f[23] = w755 ;
assign f[24] = w760 ;
assign f[25] = w765 ;
assign f[26] = w770 ;
assign f[27] = w775 ;
assign f[28] = w780 ;
assign f[29] = w785 ;
assign f[30] = w790 ;
assign f[31] = w795 ;
assign f[32] = w800 ;
assign f[33] = w805 ;
assign f[34] = w810 ;
assign f[35] = w815 ;
assign f[36] = w820 ;
assign f[37] = w825 ;
assign f[38] = w830 ;
assign f[39] = w835 ;
assign f[40] = w840 ;
assign f[41] = w845 ;
assign f[42] = w850 ;
assign f[43] = w855 ;
assign f[44] = w860 ;
assign f[45] = w865 ;
assign f[46] = w870 ;
assign f[47] = w875 ;
assign f[48] = w880 ;
assign f[49] = w885 ;
assign f[50] = w890 ;
assign f[51] = w895 ;
assign f[52] = w900 ;
assign f[53] = w905 ;
assign f[54] = w910 ;
assign f[55] = w915 ;
assign f[56] = w920 ;
assign f[57] = w925 ;
assign f[58] = w930 ;
assign f[59] = w935 ;
assign f[60] = w940 ;
assign f[61] = w945 ;
assign f[62] = w950 ;
assign f[63] = w955 ;
assign f[64] = w960 ;
assign f[65] = w965 ;
assign f[66] = w970 ;
assign f[67] = w975 ;
assign f[68] = w980 ;
assign f[69] = w985 ;
assign f[70] = w990 ;
assign f[71] = w995 ;
assign f[72] = w1000 ;
assign f[73] = w1005 ;
assign f[74] = w1010 ;
assign f[75] = w1015 ;
assign f[76] = w1020 ;
assign f[77] = w1025 ;
assign f[78] = w1030 ;
assign f[79] = w1035 ;
assign f[80] = w1040 ;
assign f[81] = w1045 ;
assign f[82] = w1050 ;
assign f[83] = w1055 ;
assign f[84] = w1060 ;
assign f[85] = w1065 ;
assign f[86] = w1070 ;
assign f[87] = w1075 ;
assign f[88] = w1080 ;
assign f[89] = w1085 ;
assign f[90] = w1090 ;
assign f[91] = w1095 ;
assign f[92] = w1100 ;
assign f[93] = w1105 ;
assign f[94] = w1110 ;
assign f[95] = w1115 ;
assign f[96] = w1120 ;
assign f[97] = w1125 ;
assign f[98] = w1130 ;
assign f[99] = w1135 ;
assign f[100] = w1140 ;
assign f[101] = w1145 ;
assign f[102] = w1150 ;
assign f[103] = w1155 ;
assign f[104] = w1160 ;
assign f[105] = w1165 ;
assign f[106] = w1170 ;
assign f[107] = w1175 ;
assign f[108] = w1180 ;
assign f[109] = w1185 ;
assign f[110] = w1190 ;
assign f[111] = w1195 ;
assign f[112] = w1200 ;
assign f[113] = w1205 ;
assign f[114] = w1210 ;
assign f[115] = w1215 ;
assign f[116] = w1220 ;
assign f[117] = w1225 ;
assign f[118] = w1230 ;
assign f[119] = w1235 ;
assign f[120] = w1240 ;
assign f[121] = w1245 ;
assign f[122] = w1250 ;
assign f[123] = w1255 ;
assign f[124] = w1260 ;
assign f[125] = w1265 ;
assign f[126] = w1270 ;
assign f[127] = w1275 ;
assign cOut = w1276 ;
endmodule
